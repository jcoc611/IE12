`timescale 1 ps / 1 ps

/**
 * Transforms an ASCII character into a 8x16 bitmap
 * of monochrome pixels.
 *
 * @param char The ASCII 7-bit character to be decoded
 * @output pixels The bitmap representing this character
 * as a 128-bit bus.
 */
module char_decoder(
	input   [`CHAR_BITES] char,
	output reg [127:0] pixels 			// TODO: should this not be FONT_BITES
);
	localparam undefined =  128'b00000000000000000000000011111111110000111010010110100101100110011001100110100101110000111111111100000000000000000000000000000000;

	always @(char) begin
		case(char)
			" ": pixels <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			"!": pixels <= undefined;
			"\"":  pixels <= undefined;
			"#":  pixels <= undefined;
			"$":  pixels <= undefined;
			"%":  pixels <= undefined;
			"&":  pixels <= undefined;
			"'":  pixels <= undefined;
			"(":  pixels <= undefined;
			")":  pixels <= undefined;
			"*":  pixels <= undefined;
			"+":  pixels <= undefined;
			",":  pixels <= undefined;
			"-":  pixels <= undefined;
			".":  pixels <= undefined;
			"/":  pixels <= undefined;
			"0":  pixels <= undefined;
			"1":  pixels <= undefined;
			"2":  pixels <= undefined;
			"3":  pixels <= undefined;
			"4":  pixels <= undefined;
			"5":  pixels <= undefined;
			"6":  pixels <= undefined;
			"7":  pixels <= undefined;
			"8":  pixels <= undefined;
			"9":  pixels <= undefined;
			":":  pixels <= undefined;
			";":  pixels <= undefined;
			"<":  pixels <= undefined;
			">":  pixels <= undefined;
			"?":  pixels <= undefined;
			"@":  pixels <= undefined;
			"A": pixels <= 128'b00000000000000000011100000111000001110000110110001101100011011000111110011000110110001101100011000000000000000000000000000000000;
			"B": pixels <= 128'b00000000000000001111110011000110110001101100011011111100110001101100011011000110110001101111110000000000000000000000000000000000;
			"C": pixels <= 128'b00000000000000000011110001100110110000001100000011000000110000001100000011000000011001100011110000000000000000000000000000000000;
			"D": pixels <= 128'b00000000000000001111100011001100110001101100011011000110110001101100011011000110110011001111100000000000000000000000000000000000;
			"E": pixels <= 128'b00000000000000001111111011000000110000001100000011111100110000001100000011000000110000001111111000000000000000000000000000000000;
			"F": pixels <= 128'b00000000000000001111111011000000110000001100000011111100110000001100000011000000110000001100000000000000000000000000000000000000;
			"G": pixels <= 128'b00000000000000000011110001100110110000001100000011000000110011101100011011000110011001100011110000000000000000000000000000000000;
			"H": pixels <= 128'b00000000000000001100011011000110110001101100011011111110110001101100011011000110110001101100011000000000000000000000000000000000;
			"I": pixels <= 128'b00000000000000000011110000011000000110000001100000011000000110000001100000011000000110000011110000000000000000000000000000000000;
			"J": pixels <= 128'b00000000000000000001111000001100000011000000110000001100000011000000110011001100110011000111100000000000000000000000000000000000;
			"K": pixels <= 128'b00000000000000001100011011001100110110001111000011100000111000001111000011011000110011001100011000000000000000000000000000000000;
			"L": pixels <= 128'b00000000000000001100000011000000110000001100000011000000110000001100000011000000110000001111111000000000000000000000000000000000;
			"M": pixels <= 128'b00000000000000001100011011101110111111101111111011010110110101101100011011000110110001101100011000000000000000000000000000000000;
			"N": pixels <= 128'b00000000000000001100011011100110111101101111111011011110110011101100011011000110110001101100011000000000000000000000000000000000;
			"O": pixels <= 128'b00000000000000000111110011000110110001101100011011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			"P": pixels <= 128'b00000000000000001111111011000110110001101100011011000110111111101100000011000000110000001100000000000000000000000000000000000000;
			"Q": pixels <= 128'b00000000000000000111110011000110110001101100011011000110110001101100011011110110110111100111110000001100000001100000000000000000;
			"R": pixels <= 128'b00000000000000001111110011000110110001101100011011000110111111001101100011001100110001101100011000000000000000000000000000000000;
			"S": pixels <= 128'b00000000000000000111110011000110110000000110000000111000000011000000011000000110110001100111110000000000000000000000000000000000;
			"T": pixels <= 128'b00000000000000000111111000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000;
			"U": pixels <= 128'b00000000000000001100011011000110110001101100011011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			"V": pixels <= 128'b00000000000000001100011011000110110001101100011001101100011011000110110000111000001110000001000000000000000000000000000000000000;
			"W": pixels <= 128'b00000000000000001100011011000110110001101100011011010110110101101111111011101110110001101100011000000000000000000000000000000000;
			"X": pixels <= 128'b00000000000000001100011011000110011011000110110000111000001110000110110001101100110001101100011000000000000000000000000000000000;
			"Y": pixels <= 128'b00000000000000000110011001100110011001100110011000111100000110000001100000011000000110000001100000000000000000000000000000000000;
			"Z": pixels <= 128'b00000000000000001111111000001100000110000001100000110000001100000110000001100000110000001111111000000000000000000000000000000000;
			"[": pixels <= undefined;
			// "\\": pixels <= undefined;
			"]": pixels <= undefined;
			"^": pixels <= undefined;
			"_": pixels <= undefined;
			"`": pixels <= undefined;
			"a": pixels <= 128'b00000000000000000000000000000000000000000111110000000110011111101100011011000110110001100111111000000000000000000000000000000000;
			"b": pixels <= 128'b00000000000000001100000011000000110000001111110011000110110001101100011011000110110001101111110000000000000000000000000000000000;
			"c": pixels <= 128'b00000000000000000000000000000000000000000111110011000110110000001100000011000000110001100111110000000000000000000000000000000000;
			"d": pixels <= 128'b00000000000000000000011000000110000001100111111011000110110001101100011011000110110001100111111000000000000000000000000000000000;
			"e": pixels <= 128'b00000000000000000000000000000000000000000111110011000110111111101100000011000000110001100111110000000000000000000000000000000000;
			"f": pixels <= 128'b00000000000000000011110001100110011000000110000011110000011000000110000001100000011000000110000000000000000000000000000000000000;
			"g": pixels <= 128'b00000000000000000000000000000000000000000111111011000110110001101100011011000110110001100111111000000110000001100111110000000000;
			"h": pixels <= 128'b00000000000000001100000011000000110000001111110011000110110001101100011011000110110001101100011000000000000000000000000000000000;
			"i": pixels <= 128'b00000000000000000001100000011000000000000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000;
			"j": pixels <= 128'b00000000000000000000011000000110000000000000011000000110000001100000011000000110000001100000011000000110011001100011110000000000;
			"k": pixels <= 128'b00000000000000001100000011000000110000001100011011001100110110001111000011011000110011001100011000000000000000000000000000000000;
			"l": pixels <= 128'b00000000000000000011100000011000000110000001100000011000000110000001100000011000000110000001100000111100000000000000000000000000;
			"m": pixels <= 128'b00000000000000000000000000000000000000001110110011010110110101101101011011010110110001101100011000000000000000000000000000000000;
			"n": pixels <= 128'b00000000000000000000000000000000000000001111110011000110110001101100011011000110110001101100011000000000000000000000000000000000;
			"o": pixels <= 128'b00000000000000000000000000000000000000000111110011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			"p": pixels <= 128'b00000000000000000000000000000000000000001111110011000110110001101100011011000110110001101111110011000000110000001100000000000000;
			"q": pixels <= 128'b00000000000000000000000000000000000000000111111011000110110001101100011011000110110001100111111000000110000001100000011000000000;
			"r": pixels <= 128'b00000000000000000000000000000000000000001111110011000110110000001100000011000000110000001100000000000000000000000000000000000000;
			"s": pixels <= 128'b00000000000000000000000000000000000000000111110011000000011100000001110000000110000001100111110000000000000000000000000000000000;
			"t": pixels <= 128'b00000000000000000001000000110000001100001111110000110000001100000011000000110000001100000001110000000000000000000000000000000000;
			"u": pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			"v": pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101100011001101100001110000001000000000000000000000000000000000000;
			"w": pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101101011011010110111111101100011000000000000000000000000000000000;
			"x": pixels <= 128'b00000000000000000000000000000000000000001100011001101100001110000011100000111000011011001100011000000000000000000000000000000000;
			"y": pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101100011011000110110001100111111000000110000001100111110000000000;
			"z": pixels <= 128'b00000000000000000000000000000000000000001111111000000110000011000001100000110000110000001111111000000000000000000000000000000000;
			"{": pixels <= undefined;
			"|": pixels <= undefined;
			"}": pixels <= undefined;
			"~": pixels <= undefined;
			default: pixels <= undefined;
		endcase
	end
endmodule
