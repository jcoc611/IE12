`timescale 1 ps / 1 ps
// Transforms an ASCII character
// into pixels (a 128 bus)
// Some Chars are not supported...

module char_decoder(
	input   [6:0] char,
	output reg [128:0] pixels
);
	localparam undefined =  128'b00000000000000000000000011111111110000111010010110100101100110011001100110100101110000111111111100000000000000000000000000000000;

	always @(char) begin
		case(char)
			// (space)
			7'b0100000: pixels <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			// !
			7'b0100001: pixels <= undefined;
			// "
			7'b0100010:  pixels <= undefined;
			// #
			7'b0100011:  pixels <= undefined;
			// $
			7'b0100100:  pixels <= undefined;
			// %
			7'b0100101:  pixels <= undefined;
			// &
			7'b0100110:  pixels <= undefined;
			// '
			7'b0100111:  pixels <= undefined;
			// (
			7'b0101000:  pixels <= undefined;
			// )
			7'b0101001:  pixels <= undefined;
			// *
			7'b0101010:  pixels <= undefined;
			// +
			7'b0101011:  pixels <= undefined;
			// ,
			7'b0101100:  pixels <= undefined;
			// -
			7'b0101101:  pixels <= undefined;
			// .
			7'b0101110:  pixels <= undefined;
			// /
			7'b0101111:  pixels <= undefined;
			// 0
			7'b0110000:  pixels <= undefined;
			// 1
			7'b0110001:  pixels <= undefined;
			// 2
			7'b0110010:  pixels <= undefined;
			// 3
			7'b0110011:  pixels <= undefined;
			// 4
			7'b0110100:  pixels <= undefined;
			// 5
			7'b0110101:  pixels <= undefined;
			// 6
			7'b0110110:  pixels <= undefined;
			// 7
			7'b0110111:  pixels <= undefined;
			// 8
			7'b0111000:  pixels <= undefined;
			// 9
			7'b0111001:  pixels <= undefined;
			// :
			7'b0111010:  pixels <= undefined;
			// ;
			7'b0111011:  pixels <= undefined;
			// <
			7'b0111100:  pixels <= undefined;
			// <=
			7'b0111101:  pixels <= undefined;
			// >
			7'b0111110:  pixels <= undefined;
			// ?
			7'b0111111:  pixels <= undefined;
			// @
			7'b1000000:  pixels <= undefined;
			// A
			7'b1000001: pixels <= 128'b00000000000000000011100000111000001110000110110001101100011011000111110011000110110001101100011000000000000000000000000000000000;
			// B
			7'b1000010: pixels <= 128'b00000000000000001111110011000110110001101100011011111100110001101100011011000110110001101111110000000000000000000000000000000000;
			// C
			7'b1000011: pixels <= 128'b00000000000000000011110001100110110000001100000011000000110000001100000011000000011001100011110000000000000000000000000000000000;
			// D
			7'b1000100: pixels <= 128'b00000000000000001111100011001100110001101100011011000110110001101100011011000110110011001111100000000000000000000000000000000000;
			// E
			7'b1000101: pixels <= 128'b00000000000000001111111011000000110000001100000011111100110000001100000011000000110000001111111000000000000000000000000000000000;
			// F
			7'b1000110: pixels <= 128'b00000000000000001111111011000000110000001100000011111100110000001100000011000000110000001100000000000000000000000000000000000000;
			// G
			7'b1000111: pixels <= 128'b00000000000000000011110001100110110000001100000011000000110011101100011011000110011001100011110000000000000000000000000000000000;
			// H
			7'b1001000: pixels <= 128'b00000000000000001100011011000110110001101100011011111110110001101100011011000110110001101100011000000000000000000000000000000000;
			// I
			7'b1001001: pixels <= 128'b00000000000000000011110000011000000110000001100000011000000110000001100000011000000110000011110000000000000000000000000000000000;
			// J
			7'b1001010: pixels <= 128'b00000000000000000001111000001100000011000000110000001100000011000000110011001100110011000111100000000000000000000000000000000000;
			// K
			7'b1001011: pixels <= 128'b00000000000000001100011011001100110110001111000011100000111000001111000011011000110011001100011000000000000000000000000000000000;
			// L
			7'b1001100: pixels <= 128'b00000000000000001100000011000000110000001100000011000000110000001100000011000000110000001111111000000000000000000000000000000000;
			// M
			7'b1001101: pixels <= 128'b00000000000000001100011011101110111111101111111011010110110101101100011011000110110001101100011000000000000000000000000000000000;
			// N
			7'b1001110: pixels <= 128'b00000000000000001100011011100110111101101111111011011110110011101100011011000110110001101100011000000000000000000000000000000000;
			// O
			7'b1001111: pixels <= 128'b00000000000000000111110011000110110001101100011011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			// P
			7'b1010000: pixels <= 128'b00000000000000001111111011000110110001101100011011000110111111101100000011000000110000001100000000000000000000000000000000000000;
			// Q
			7'b1010001: pixels <= 128'b00000000000000000111110011000110110001101100011011000110110001101100011011110110110111100111110000001100000001100000000000000000;
			// R
			7'b1010010: pixels <= 128'b00000000000000001111110011000110110001101100011011000110111111001101100011001100110001101100011000000000000000000000000000000000;
			// S
			7'b1010011: pixels <= 128'b00000000000000000111110011000110110000000110000000111000000011000000011000000110110001100111110000000000000000000000000000000000;
			// T
			7'b1010100: pixels <= 128'b00000000000000000111111000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000;
			// U
			7'b1010101: pixels <= 128'b00000000000000001100011011000110110001101100011011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			// V
			7'b1010110: pixels <= 128'b00000000000000001100011011000110110001101100011001101100011011000110110000111000001110000001000000000000000000000000000000000000;
			// W
			7'b1010111: pixels <= 128'b00000000000000001100011011000110110001101100011011010110110101101111111011101110110001101100011000000000000000000000000000000000;
			// X
			7'b1011000: pixels <= 128'b00000000000000001100011011000110011011000110110000111000001110000110110001101100110001101100011000000000000000000000000000000000;
			// Y
			7'b1011001: pixels <= 128'b00000000000000000110011001100110011001100110011000111100000110000001100000011000000110000001100000000000000000000000000000000000;
			// Z
			7'b1011010: pixels <= 128'b00000000000000001111111000001100000110000001100000110000001100000110000001100000110000001111111000000000000000000000000000000000;
			// [
			7'b1011011: pixels <= undefined;
			// \
			7'b1011100: pixels <= undefined;
			// ]
			7'b1011101: pixels <= undefined;
			// ^
			7'b1011110: pixels <= undefined;
			// _
			7'b1011111: pixels <= undefined;
			// `
			7'b1100000: pixels <= undefined;
			// a
			7'b1100001: pixels <= 128'b00000000000000000000000000000000000000000111110000000110011111101100011011000110110001100111111000000000000000000000000000000000;
			// b
			7'b1100010: pixels <= 128'b00000000000000001100000011000000110000001111110011000110110001101100011011000110110001101111110000000000000000000000000000000000;
			// c
			7'b1100011: pixels <= 128'b00000000000000000000000000000000000000000111110011000110110000001100000011000000110001100111110000000000000000000000000000000000;
			 // d
			7'b1100100: pixels <= 128'b00000000000000000000011000000110000001100111111011000110110001101100011011000110110001100111111000000000000000000000000000000000;
			 // e
			7'b1100101: pixels <= 128'b00000000000000000000000000000000000000000111110011000110111111101100000011000000110001100111110000000000000000000000000000000000;
			 // f
			7'b1100110: pixels <= 128'b00000000000000000011110001100110011000000110000011110000011000000110000001100000011000000110000000000000000000000000000000000000;
			 // g
			7'b1100111: pixels <= 128'b00000000000000000000000000000000000000000111111011000110110001101100011011000110110001100111111000000110000001100111110000000000;
			// h
			7'b1101000: pixels <= 128'b00000000000000001100000011000000110000001111110011000110110001101100011011000110110001101100011000000000000000000000000000000000;
			 // i
			7'b1101001: pixels <= 128'b00000000000000000001100000011000000000000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000;
			 // j
			7'b1101010: pixels <= 128'b00000000000000000000011000000110000000000000011000000110000001100000011000000110000001100000011000000110011001100011110000000000;
			 // k
			7'b1101011: pixels <= 128'b00000000000000001100000011000000110000001100011011001100110110001111000011011000110011001100011000000000000000000000000000000000;
			 // l
			7'b1101100: pixels <= 128'b00000000000000000011100000011000000110000001100000011000000110000001100000011000000110000001100000111100000000000000000000000000;
			 // m
			7'b1101101: pixels <= 128'b00000000000000000000000000000000000000001110110011010110110101101101011011010110110001101100011000000000000000000000000000000000;
			 // n
			7'b1101110: pixels <= 128'b00000000000000000000000000000000000000001111110011000110110001101100011011000110110001101100011000000000000000000000000000000000;
			 // o
			7'b1101111: pixels <= 128'b00000000000000000000000000000000000000000111110011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			 // p
			7'b1110000: pixels <= 128'b00000000000000000000000000000000000000001111110011000110110001101100011011000110110001101111110011000000110000001100000000000000;
			// q
			7'b1110001: pixels <= 128'b00000000000000000000000000000000000000000111111011000110110001101100011011000110110001100111111000000110000001100000011000000000;
			 // r
			7'b1110010: pixels <= 128'b00000000000000000000000000000000000000001111110011000110110000001100000011000000110000001100000000000000000000000000000000000000;
			 // s
			7'b1110011: pixels <= 128'b00000000000000000000000000000000000000000111110011000000011100000001110000000110000001100111110000000000000000000000000000000000;
			 // t
			7'b1110100: pixels <= 128'b00000000000000000001000000110000001100001111110000110000001100000011000000110000001100000001110000000000000000000000000000000000;
			 // u
			7'b1110101: pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101100011011000110110001100111110000000000000000000000000000000000;
			 // v
			7'b1110110: pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101100011001101100001110000001000000000000000000000000000000000000;
			 // w
			7'b1110111: pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101101011011010110111111101100011000000000000000000000000000000000;
			 // x
			7'b1111000: pixels <= 128'b00000000000000000000000000000000000000001100011001101100001110000011100000111000011011001100011000000000000000000000000000000000;
			 // y
			7'b1111001: pixels <= 128'b00000000000000000000000000000000000000001100011011000110110001101100011011000110110001100111111000000110000001100111110000000000;
			 // z
			7'b1111010: pixels <= 128'b00000000000000000000000000000000000000001111111000000110000011000001100000110000110000001111111000000000000000000000000000000000;
			 // {
			7'b1111011: pixels <= undefined;
			 // |
			7'b1111100: pixels <= undefined;
			 // }
			7'b1111101: pixels <= undefined;
			 // ~
			7'b1111110: pixels <= undefined;
			default: pixels <= undefined;
		endcase
	end
endmodule
